`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.09.2016 08:48:06
// Design Name: 
// Module Name: manager
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ipManager(
    // implementation of AXI Slave interface
    /*input S00_AXI_awaddr,
    input S00_AXI_awlen, 
    input S00_AXI_awsize,
    input S00_AXI_awburst,
    input S00_AXI_awlock,
    input S00_AXI_awcache,
    input S00_AXI_awprot,
    input S00_AXI_awregion,
    input S00_AXI_awqos,
    input S00_AXI_awvalid,
    output S00_AXI_awready,
    input S00_AXI_awdata,
    input S00_AXI_awstrb,
    input S00_AXI_awlast,
    input S00_AXI_wvalid,
    output S00_AXI_awready,
    output S00_AXI_bresp,
    output S00_AXI_bvalid,
    input S00_AXI_bready,
    input S00_AXI_arradr,
    input S00_AXI_arlen,
    input S00_AXI_arsize,
    input S00_AXI_arburst,
    input S00_AXI_arlock,
    input S00_AXI_arcache,
    input S00_AXI_arprot,
    input S00_AXI_arregion,
    input S00_AXI_arqos,
    input S00_AXI_arvalid,
    output S00_AXI_arready,
    output S00_AXI_rdata,
    output S00_AXI_rresp,
    output S00_AXI_rlast,
    output S00_AXI_rvalid,
    input S00_AXI_rready,*/
    // custom logic
    output enable
    );
endmodule
